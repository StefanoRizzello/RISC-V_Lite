-------------------------------------------------------------------------------
-- Title      : unary_AND
-- Project    : 
-------------------------------------------------------------------------------
-- File       : unary_AND.vhd
-- Author     : GR17 (F.Bongo, S.Rizzello, F.Vacca)
-- Company    : 
-- Created    : 2022-01-21
-- Last update: 2022-02-01
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2022 
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

-------------------------------------------------------------------------------

entity unary_AND is

  port (
    inp  : in  std_logic_vector(31 downto 0);
    outp : out std_logic);

end entity unary_AND;

-------------------------------------------------------------------------------

architecture str of unary_AND is

  -----------------------------------------------------------------------------
  -- Internal signal declarations
  -----------------------------------------------------------------------------

  signal temp : std_logic_vector(31 downto 0);

begin  -- architecture str

  temp(0) <= inp(0);
  gen : for i in 1 to 31 generate
          temp(i) <= temp(i-1) and inp(i);
        end generate;
  outp <= temp(31);

  -----------------------------------------------------------------------------
  -- Component instantiations
  -----------------------------------------------------------------------------

end architecture str;

-------------------------------------------------------------------------------
